module freq_divider();
	input
	output
	
endmodule 